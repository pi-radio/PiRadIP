package piradma_mm2s;

endpackage